`ifndef SLAVE_AGENT_BFM_INCLUDED_
`define SLAVE_AGENT_BFM_INCLUDED_

//--------------------------------------------------------------------------------------------
// Module : Slave Agent BFM 
// This module is used as the configuration class for slave agent bfm and its components
//--------------------------------------------------------------------------------------------
module slave_agent_bfm(spi_if intf);

  //-------------------------------------------------------
  // Package : Importing Uvm Pakckage and Test Package
  //-------------------------------------------------------
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //-------------------------------------------------------
  // Slave driver bfm instantiation
  //-------------------------------------------------------
  //slave_driver_bfm slave_drv_bfm_h (.sclk(intf.sclk),.cs(intf.cs),.mosi(intf.mosi),.miso(intf.miso));
  slave_driver_bfm slave_drv_bfm_h (intf);

 //-------------------------------------------------------
  // Slave monitor bfm instantiation
  //-------------------------------------------------------
  //slave_monitor_bfm slave_mon_bfm_h (.sclk(intf.sclk),.mosi(intf.miso));
  slave_monitor_bfm slave_mon_bfm_h (intf);

  //-------------------------------------------------------
  // Setting Slave_driver_bfm and monitor_bfm
  //-------------------------------------------------------
  initial begin
    uvm_config_db#(virtual slave_driver_bfm)::set(null,"*", "slave_driver_bfm", slave_drv_bfm_h); 
    uvm_config_db#(virtual slave_monitor_bfm)::set(null,"*", "slave_monitor_bfm", slave_mon_bfm_h); 
  end

  initial begin
    $display("Slave Agent BFM");
  end

endmodule : slave_agent_bfm

`endif
