//-------------------------------------------------------
//Here declaring the interface as spi_if
//-------------------------------------------------------


  interface spi_if;

    logic sclock;
    logic mosi;
    logic miso;
    logic ss;

    //-------------------------------------------------------
    //Here we are declaring clocking block and mod modports
    //-------------------------------------------------------

  endinterface
