//-------------------------------------------------------
//
//top
//-------------------------------------------------------
