In this test we are starting the spi_fd_8b_vseq on the virtula sequencer
