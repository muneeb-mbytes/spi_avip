`define SIZE 3
`define DW 2**`SIZE
