module master_drv;

virtual spi_if vif;




endmodule
