 module master_agent_bfm

 `include master_drv drv_h(in1);
 `include master_mon mon_h(in1);




 endmodule
