Testing if the lock works on phase1_development_branch
