Testing to see if main lock is enabled
