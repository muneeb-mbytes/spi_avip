`ifndef SPI_FD_CONFIG_CPOL1_CPHA1_MSB_C2T_T2C_BAUDRATE_MASTER_SEQ_INCLUDED_
`define SPI_FD_CONFIG_CPOL1_CPHA1_MSB_C2T_T2C_BAUDRATE_MASTER_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// class: extended class from base class
//--------------------------------------------------------------------------------------------
class spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq extends master_base_seq;

  //register with factory so can use create uvm_method 
  //and override in future if necessary 

   `uvm_object_utils(spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq)

  //---------------------------------------------
  // Externally defined tasks and functions
  //---------------------------------------------

   extern function new (string name="spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq");

   extern virtual task body();
endclass:spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq

//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_sequence class object
//
// Parameters:
//  name - instance name of the config_template
//-----------------------------------------------------------------------------
function spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq::new(string name="spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq");
  super.new(name);
endfunction:new

//-----------------------------------------------------------------------------
//task:body
//based on the request from driver task will drive the transaction
//-----------------------------------------------------------------------------
task spi_fd_config_cpol1_cpha1_msb_c2t_t2c_baudrate_master_seq::body(); 
  req=master_tx::type_id::create("req");
  start_item(req);
  if(!req.randomize() with {req.master_out_slave_in.size() == 1;
                            // selecting only one slave  
                            $countones(req.cs) == NO_OF_SLAVES - 1;
                            // selecting slave 0
                            req.cs[0] == 0;
                           }) begin
    `uvm_fatal(get_type_name(),"Randomization failed")
  end
  `uvm_info(get_type_name(),$sformatf("master_seq",req.sprint()),UVM_MEDIUM)
  finish_item(req);

endtask:body

`endif

