//--------------------------------------------------------------------------------------------
// Module       : Slave Driver BFM
// Description  : Connects the slave driver bfm with the driver proxy
//--------------------------------------------------------------------------------------------
module slave_driver_bfm(spi_if intf);

  initial begin
    $display("Slave Driver BFM");
  end

endmodule : slave_driver_bfm
