Testing if the lock works on phase1_development_branch
Adding changes to see at Chetan's workspace area 
