//-------------------------------------------------------
//master monitor
//-------------------------------------------------------
module master_mon(spi_intf);

  initial
  begin
    $display("Master Monitor BFM");
  end

endmodule
