module master_mon;

virtual spi_if vif;


endmodule
