`ifndef SPI_QUAD_SPI_TYPE_VIRTUAL_SEQ_INCLUDED_
`define SPI_QUAD_SPI_TYPE_VIRTUAL_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Extended class from spi virtual sequence
//--------------------------------------------------------------------------------------------
class spi_quad_spi_type_virtual_seq extends spi_fd_virtual_seq_base;
  
  `uvm_object_utils(spi_quad_spi_type_virtual_seq)

  //declare extended class handles of master and slave sequence
  spi_quad_spi_type_master_seq spi_quad_spi_type_master_seq_h;
  spi_quad_spi_type_slave_seq spi_quad_spi_type_slave_seq_h;

  //--------------------------------------------------------------------------------------------
  // Externally defined tasks and functions
  //--------------------------------------------------------------------------------------------
  extern function new(string name="spi_quad_spi_type_virtual_seq");
  extern task body();

endclass : spi_quad_spi_type_virtual_seq

//--------------------------------------------------------------------------------------------
//Constructor:new
//
//Paramters:
//name - Instance name of the virtual_sequence
//parent - parent under which this component is created
//--------------------------------------------------------------------------------------------
function spi_quad_spi_type_virtual_seq::new(string name="spi_quad_spi_type_virtual_seq");
  super.new(name);
endfunction: new

//--------------------------------------------------------------------------------------------
//task:body
//Creates the required ports
//
//Parameters:
// phase - stores the current phase
//--------------------------------------------------------------------------------------------
task spi_quad_spi_type_virtual_seq::body();
 super.body(); //Sets up the sub-sequencer pointer
 
 //crearions master and slave sequence handles here  
 spi_quad_spi_type_master_seq_h=spi_quad_spi_type_master_seq::type_id::create("spi_quad_spi_type_master_seq_h");
 spi_quad_spi_type_slave_seq_h=spi_quad_spi_type_slave_seq::type_id::create("spi_quad_spi_type_slave_seq_h");

    //configuring no of masters and starting master sequencers

  fork
     // TODO(mshariff): We need to connect the slaves with caution
      // as only ONe slave can drive on MISO line
      // so the sequences need to be started based on the System configurations

      // MSHA: //has_s_agt should be declared in env_config file
      // MSHA: if(e_cfg_h.has_s_agt) begin 
      // MSHA:   //no_of_sagent should be declared in env_config file
      // MSHA: for(int i=0; i<e_cfg_h.no_of_sagent; i++)begin
      // MSHA:   //starting slave sequencer
      // MSHA:  spi_quad_spi_type_slave_seq_h.start(s_seqr_h);
      // MSHA:  end
      // MSHA: end

      //starting slave sequencer
      forever begin: SLAVE_SEQ_START
        spi_quad_spi_type_slave_seq_h.start(p_sequencer.slave_seqr_h);
      end
    join_none
    //has_m_agt should be declared in env_config file
    // TODO(mshariff): Only one Master agent as SPI supports only one Master

    // MSHA: if(e_cfg_h.has_m_agt)begin
    // MSHA: //no_of_magent should be declared in env_config file
    // MSHA: for(int i=0; i<e_cfg_h.no_of_magent; i++)begin
    // MSHA:   //starting master sequencer
    // MSHA:   spi_quad_spi_type_master_seq_h.start(m_seqr_h);
    // MSHA:   end
    // MSHA: end

    //starting master sequencer
    repeat(5)begin: MASTER_SEQ_START
      spi_quad_spi_type_master_seq_h.start(p_sequencer.master_seqr_h);
    end

endtask: body

`endif
